package pds_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   
   `include "coverage.svh"
   `include "base_tester.svh"
   `include "random_tester.svh"
   `include "cpwr_tester.svh"   
   `include "scoreboard.svh"
   `include "env.svh"
   `include "random_test.svh"
   `include "cpwr_test.svh"
   
endpackage : pds_pkg
